library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity clk_div is
    Port (  
        clk : in std_logic;
        sclk : out std_logic
    );
end clk_div;

architecture my_clk_div of clk_div is
    constant max_count : integer := (1100);    
    signal tmp_clk : std_logic := '0';
begin
    my_div: process (clk)
        variable div_cnt : integer := 0;
    begin
        if (rising_edge(clk)) then
            if (div_cnt = MAX_COUNT) then
                tmp_clk <= not tmp_clk;
                div_cnt := 0;
            else
                div_cnt := div_cnt + 1;
            end if;
        end if;
    end process my_div;
    
    sclk <= tmp_clk;
end my_clk_div;
